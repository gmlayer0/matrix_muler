`timescale 1ps/1ps

module axi_raw_bram_wrap #(
    parameter int bram_size = ,
    parameter  = ,
)(
    input clk,
    input rst,

);
    
endmodule